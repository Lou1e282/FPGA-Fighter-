module player_jump #(

)
(

); 

endmodule