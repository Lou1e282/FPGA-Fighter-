module player_hp (
    
    

)


endmodule